module Binary_to_BCD
(
	input wire [15:0] binary,
	output wire [15:0] BCD_code
);
//jdsklfjskl
wire [3:0] a1,a2,a3,a4,a5,a6,a7;
wire [3:0] b1,b2,b3,b4,b5,b6,b7;

assign b1 = {1'b0,binary[7:5]};
assign b2 = {a1[2:0],binary[4]};
assign b3 = {a2[2:0],binary[3]};
assign b4 = {a3[2:0],binary[2]};
assign b5 = {a4[2:0],binary[1]};
assign b6 = {1'b0,a1[3],a2[3],a3[3]};
assign b7 = {a6[2:0],a4[3]};

assign a1 = b1 == 4'b0101 ? 4'b1000 : (b1 == 4'b0110 ? 4'b1001 : (b1 == 4'b0111 ? 4'b1010 : (b1 == 4'b1000 ? 4'b1011 : b1 == 4'b1001 ? 4'b1100 : b1)));
assign a2 = b2 == 4'b0101 ? 4'b1000 : (b2 == 4'b0110 ? 4'b1001 : (b2 == 4'b0111 ? 4'b1010 : (b2 == 4'b1000 ? 4'b1011 : b2 == 4'b1001 ? 4'b1100 : b2)));
assign a3 = b3 == 4'b0101 ? 4'b1000 : (b3 == 4'b0110 ? 4'b1001 : (b3 == 4'b0111 ? 4'b1010 : (b3 == 4'b1000 ? 4'b1011 : b3 == 4'b1001 ? 4'b1100 : b3)));
assign a4 = b4 == 4'b0101 ? 4'b1000 : (b4 == 4'b0110 ? 4'b1001 : (b4 == 4'b0111 ? 4'b1010 : (b4 == 4'b1000 ? 4'b1011 : b4 == 4'b1001 ? 4'b1100 : b4)));
assign a5 = b5 == 4'b0101 ? 4'b1000 : (b5 == 4'b0110 ? 4'b1001 : (b5 == 4'b0111 ? 4'b1010 : (b5 == 4'b1000 ? 4'b1011 : b5 == 4'b1001 ? 4'b1100 : b5)));
assign a6 = b6 == 4'b0101 ? 4'b1000 : (b6 == 4'b0110 ? 4'b1001 : (b6 == 4'b0111 ? 4'b1010 : (b6 == 4'b1000 ? 4'b1011 : b6 == 4'b1001 ? 4'b1100 : b6)));
assign a7 = b7 == 4'b0101 ? 4'b1000 : (b7 == 4'b0110 ? 4'b1001 : (b7 == 4'b0111 ? 4'b1010 : (b7 == 4'b1000 ? 4'b1011 : b7 == 4'b1001 ? 4'b1100 : b7)));

assign BCD_code = {2'd0,a6[3],a7[3],a7[2:0],a5[3],a5[2:0],binary[0],4'd0};

endmodule
